module not_gate (
    input logic a,    // Вход a
    output logic y    // Выход y
);
    assign y = ~a;    // Логическая операция NOT
endmodule
